// Level 10 - Advanced Logic Design
// TODO: Implement a complex multiplexer
// This is an editable file for level 10

module advanced_mux (
    input [3:0] data,
    input [1:0] sel,
    output y
);
    // Your implementation here
    
endmodule