// Level 1 - Basic Gate Implementation
// TODO: Implement a simple AND gate
// Inputs: a, b
// Output: y

module and_gate (
    input a,
    input b,
    output y
);
    // Your implementation here
    
endmodule